/*-------------------------------------------------------------------------
// Module:  rom
// File:    rom.sv
// Author:  shawn Liu
// E-mail:  shawn110285@gmail.com
// Description: two ports rom, one port for lsu read and the other for instruction
//              fetch
--------------------------------------------------------------------------*/

// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------

//`include "../../core/include/defines.v"
`include "defines.v"

module rom(
	input wire				      rom_clk_i,
    input wire                    rom_n_rst_i,
	input wire					  rom_ce_i,
	input wire[`DataAddrBus]	  rom_addr_i,
	output reg[`DataBus]		  rom_data_o,

    // lsu data port
	input wire				      clk_i,
	input wire                    n_rst_i,
	input wire					  ce_i,
	input wire[3:0]				  sel_i,
	input wire[`DataAddrBus]	  addr_i,
	input wire					  we_i,
	input wire[`DataBus]		  data_i,
	output wire                   rvalid_o,
	output reg[`DataBus]		  data_o
);

    /* verilator lint_off LITENDIAN */
    logic [0:`RomNum-1][`InstBus]  rom_mem;
    /* verilator lint_on LITENDIAN */

    assign rvalid_o = ce_i & (~we_i);
    // the content is from the boot rom
    assign rom_mem =
    {
     32'h3050006f,
     32'h3010006f,
     32'h2fd0006f,
     32'h2f90006f,
     32'h2f50006f,
     32'h2f10006f,
     32'h2ed0006f,
     32'h2e90006f,
     32'h2e50006f,
     32'h2e10006f,
     32'h2dd0006f,
     32'h2d90006f,
     32'h2d50006f,
     32'h2d10006f,
     32'h2cd0006f,
     32'h2c90006f,
     32'h2c50006f,
     32'h2c10006f,
     32'h2bd0006f,
     32'h2b90006f,
     32'h2b50006f,
     32'h2b10006f,
     32'h2ad0006f,
     32'h2a90006f,
     32'h2a50006f,
     32'h2a10006f,
     32'h29d0006f,
     32'h2990006f,
     32'h2950006f,
     32'h2910006f,
     32'h28d0006f,
     32'h2890006f,
     32'h3990006f,
     32'h000057b7,
     32'h1b800713,
     32'h00e7a423,
     32'h00300713,
     32'h00e7a023,
     32'h00008067,
     32'h00005737,
     32'h00472783,
     32'h0017f793,
     32'hfe079ce3,
     32'h000057b7,
     32'h00a7a623,
     32'h00008067,
     32'hff010113,
     32'h00112623,
     32'h00812423,
     32'h00912223,
     32'h01212023,
     32'h00050493,
     32'h00800413,
     32'h00900913,
     32'h0180006f,
     32'h03750513,
     32'hfbdff0ef,
     32'h00449493,
     32'hfff40413,
     32'h00040c63,
     32'h01c4d513,
     32'hfea944e3,
     32'h03050513,
     32'hfa1ff0ef,
     32'hfe5ff06f,
     32'h00c12083,
     32'h00812403,
     32'h00412483,
     32'h00012903,
     32'h01010113,
     32'h00008067,
     32'hff010113,
     32'h00112623,
     32'h00812423,
     32'h00050413,
     32'h00054503,
     32'h00050a63,
     32'hf69ff0ef,
     32'h00140413,
     32'h00044503,
     32'hfe051ae3,
     32'h00c12083,
     32'h00812403,
     32'h01010113,
     32'h00008067,
     32'h000057b7,
     32'h0047a503,
     32'h00257513,
     32'h00008067,
     32'h00005737,
     32'h00472783,
     32'h0027f793,
     32'hfe078ce3,
     32'h000057b7,
     32'h0007a223,
     32'h0107a503,
     32'h0ff57513,
     32'h00008067,
     32'hfe010113,
     32'h00112e23,
     32'h00812c23,
     32'h00912a23,
     32'h01212823,
     32'h01312623,
     32'h01412423,
     32'h00050a13,
     32'h00058993,
     32'h00000413,
     32'h00d00493,
     32'h00a00913,
     32'hfadff0ef,
     32'h00950e63,
     32'h01250c63,
     32'hff347ae3,
     32'h008a07b3,
     32'h00a78023,
     32'h00140413,
     32'hfe5ff06f,
     32'h00a00513,
     32'hec1ff0ef,
     32'h008a0433,
     32'h00040023,
     32'h01c12083,
     32'h01812403,
     32'h01412483,
     32'h01012903,
     32'h00c12983,
     32'h00812a03,
     32'h02010113,
     32'h00008067,
     32'h00002717,
     32'hdf870713,
     32'h00072783,
     32'h00178793,
     32'h00f72023,
     32'h00008067,
     32'hfc010113,
     32'h02112e23,
     32'h02812c23,
     32'h02912a23,
     32'h03212823,
     32'h03312623,
     32'h03412423,
     32'h03512223,
     32'h03612023,
     32'h01712e23,
     32'h01812c23,
     32'h00012423,
     32'h00010623,
     32'h00006437,
     32'h00400793,
     32'h00f42223,
     32'he25ff0ef,
     32'h00800793,
     32'h00f42223,
     32'h00001797,
     32'hd7c78793,
     32'h0007a503,
     32'hea5ff0ef,
     32'h00300793,
     32'h00f42223,
     32'h250000ef,
     32'h00600793,
     32'h00f42223,
     32'h00000617,
     32'hf7860613,
     32'h02faf537,
     32'h08050513,
     32'h00000593,
     32'h388000ef,
     32'h00700793,
     32'h00f42223,
     32'h00002797,
     32'hd4078c23,
     32'h00002797,
     32'hd407a423,
     32'h00002417,
     32'hd4840413,
     32'h00001a17,
     32'hd24a0a13,
     32'h00001917,
     32'hd2090913,
     32'h00001497,
     32'ha1448493,
     32'h07300993,
     32'h00001a97,
     32'hb40a8a93,
     32'h00044783,
     32'h00100613,
     32'h01879693,
     32'h4186d693,
     32'h00400713,
     32'h08c78c63,
     32'h02068863,
     32'hfee79ce3,
     32'h000067b7,
     32'h00200713,
     32'h00e7a223,
     32'h00001517,
     32'hb5050513,
     32'hdfdff0ef,
     32'h00001517,
     32'hb7050513,
     32'hdf1ff0ef,
     32'h0000006f,
     32'h00002797,
     32'hccc78793,
     32'h0007a783,
     32'h00500713,
     32'h00f77863,
     32'h00400793,
     32'h00f40023,
     32'hf9dff06f,
     32'h00600593,
     32'h40f585b3,
     32'h00001517,
     32'haac50513,
     32'h764000ef,
     32'hdedff0ef,
     32'hf80500e3,
     32'hdf5ff0ef,
     32'h00100793,
     32'h00f40023,
     32'h00001797,
     32'hc7878793,
     32'h0007a503,
     32'hd95ff0ef,
     32'h00092503,
     32'hd8dff0ef,
     32'hf59ff06f,
     32'h00500593,
     32'h00810513,
     32'hde9ff0ef,
     32'h00810513,
     32'hd75ff0ef,
     32'h00914783,
     32'h02079663,
     32'h00814783,
     32'hfbc78793,
     32'h0ff7f693,
     32'h02f00713,
     32'h0ed76e63,
     32'h00269793,
     32'h009787b3,
     32'h0007a783,
     32'h009787b3,
     32'h00078067,
     32'h000a2503,
     32'hd3dff0ef,
     32'h00092503,
     32'hd35ff0ef,
     32'h00810b13,
     32'h00d10c13,
     32'h00001b97,
     32'ha44b8b93,
     32'h000b4503,
     32'hc9dff0ef,
     32'h000b8513,
     32'hd15ff0ef,
     32'h001b0b13,
     32'hff6c16e3,
     32'hed9ff06f,
     32'h06e00513,
     32'hc81ff0ef,
     32'h06600c13,
     32'hd41ff0ef,
     32'h03850863,
     32'h05351063,
     32'hd35ff0ef,
     32'h00050b93,
     32'h00050a63,
     32'h00000b13,
     32'hd25ff0ef,
     32'h001b0b13,
     32'hff7b1ce3,
     32'h06e00513,
     32'hc4dff0ef,
     32'hfd1ff06f,
     32'h06e00513,
     32'hc41ff0ef,
     32'h00092503,
     32'hcb9ff0ef,
     32'he85ff06f,
     32'h000a8513,
     32'hcadff0ef,
     32'hfb1ff06f,
     32'h00092503,
     32'hca1ff0ef,
     32'h00001517,
     32'h9bc50513,
     32'hc95ff0ef,
     32'h00000513,
     32'h048000ef,
     32'h02e00513,
     32'hc05ff0ef,
     32'h00001517,
     32'h9b850513,
     32'hc79ff0ef,
     32'h00092503,
     32'hc71ff0ef,
     32'he3dff06f,
     32'h00400793,
     32'h00f40023,
     32'he31ff06f,
     32'h000a2503,
     32'hc59ff0ef,
     32'h00092503,
     32'hc51ff0ef,
     32'he1dff06f,
     32'h00008067,
     32'h00008067,
     32'h00008067,
     32'hff010113,
     32'h00112623,
     32'h0f0000ef,
     32'h00f57513,
     32'h000067b7,
     32'h00a7a223,
     32'h00001517,
     32'ha7050513,
     32'hc1dff0ef,
     32'h00001517,
     32'ha7c50513,
     32'hc11ff0ef,
     32'h00001517,
     32'ha8050513,
     32'hc05ff0ef,
     32'h0cc000ef,
     32'hb99ff0ef,
     32'h00001517,
     32'ha7c50513,
     32'hbf1ff0ef,
     32'h0a0000ef,
     32'hb85ff0ef,
     32'h00001517,
     32'ha7850513,
     32'hbddff0ef,
     32'h094000ef,
     32'hb71ff0ef,
     32'h00001517,
     32'ha7450513,
     32'hbc9ff0ef,
     32'h088000ef,
     32'hb5dff0ef,
     32'h00001517,
     32'ha7050513,
     32'hbb5ff0ef,
     32'h0000006f,
     32'hff010113,
     32'h00112623,
     32'h00812423,
     32'h342026f3,
     32'h800007b7,
     32'h00778793,
     32'h04d79263,
     32'h000067b7,
     32'h0007a403,
     32'h110000ef,
     32'h00447793,
     32'h02078063,
     32'hffb47413,
     32'h000067b7,
     32'h0087a223,
     32'h00c12083,
     32'h00812403,
     32'h01010113,
     32'h00008067,
     32'h00446413,
     32'h000067b7,
     32'h0087a223,
     32'hfe5ff06f,
     32'hf15ff0ef,
     32'h34102573,
     32'h00008067,
     32'h34202573,
     32'h00008067,
     32'h34302573,
     32'h00008067,
     32'h30502573,
     32'h00008067,
     32'hc0002573,
     32'hc80025f3,
     32'h00008067,
     32'h000047b7,
     32'h0047a583,
     32'h0007a503,
     32'h0047a703,
     32'hfeb71ae3,
     32'h00008067,
     32'h000047b7,
     32'hfff00713,
     32'h00e7a423,
     32'h00b7a623,
     32'h00a7a423,
     32'h00008067,
     32'hff010113,
     32'h00112623,
     32'h00812423,
     32'h00912223,
     32'h00050413,
     32'h00058493,
     32'h000067b7,
     32'h00f00713,
     32'h00e7a223,
     32'h00002797,
     32'h9c078793,
     32'h00a7a023,
     32'h00b7a223,
     32'h00002797,
     32'h9ac7a223,
     32'hf95ff0ef,
     32'h00a40533,
     32'h00853433,
     32'h00b485b3,
     32'h00b405b3,
     32'hf99ff0ef,
     32'h08000793,
     32'h3047a073,
     32'h00800793,
     32'h3007a073,
     32'h00c12083,
     32'h00812403,
     32'h00412483,
     32'h01010113,
     32'h00008067,
     32'hff010113,
     32'h00112623,
     32'h00812423,
     32'h00912223,
     32'h00002797,
     32'h95c78793,
     32'h0007a403,
     32'h0047a483,
     32'hf39ff0ef,
     32'h00a40533,
     32'h00853433,
     32'h00b485b3,
     32'h00b405b3,
     32'hf3dff0ef,
     32'h00002797,
     32'h92878793,
     32'h0007a783,
     32'h00078463,
     32'h000780e7,
     32'h00c12083,
     32'h00812403,
     32'h00412483,
     32'h01010113,
     32'h00008067,
     32'h08000793,
     32'h3047b073,
     32'h00008067,
     32'hfb010113,
     32'h04112623,
     32'h04812423,
     32'h04912223,
     32'h05212023,
     32'h03312e23,
     32'h03412c23,
     32'h03512a23,
     32'h03612823,
     32'h03712623,
     32'h03812423,
     32'h03912223,
     32'h03a12023,
     32'h01b12e23,
     32'h00050413,
     32'h00058a13,
     32'h02500a93,
     32'h03000b93,
     32'h00900493,
     32'h00000b17,
     32'h650b0b13,
     32'h01000993,
     32'h00010913,
     32'h00c0006f,
     32'h00140413,
     32'h929ff0ef,
     32'h00044503,
     32'h30050863,
     32'hff5518e3,
     32'h00144503,
     32'h09750a63,
     32'h02d00793,
     32'h08f50e63,
     32'h00240413,
     32'h00000813,
     32'hfd050793,
     32'h0ff7f793,
     32'h08f4ec63,
     32'h00000c93,
     32'h002c9793,
     32'h019787b3,
     32'h00179793,
     32'h00a787b3,
     32'hfd078c93,
     32'h00140413,
     32'hfff44503,
     32'hfd050793,
     32'h0ff7f793,
     32'hfcf4fee3,
     32'h0df57793,
     32'h04c00713,
     32'h06e78463,
     32'h2a050663,
     32'h06000793,
     32'h00050613,
     32'h00a7f663,
     32'hfe050613,
     32'h0ff67613,
     32'hfbe60793,
     32'h0ff7f693,
     32'h01600713,
     32'h0ed76a63,
     32'h00269793,
     32'h016787b3,
     32'h0007a783,
     32'h016787b3,
     32'h00078067,
     32'h00244503,
     32'h00340413,
     32'h00100813,
     32'hf75ff06f,
     32'h00244503,
     32'h00340413,
     32'h00200813,
     32'hf65ff06f,
     32'h00000c93,
     32'hf95ff06f,
     32'h00486813,
     32'h00044503,
     32'h00140413,
     32'hf91ff06f,
     32'h004a0c13,
     32'h000a2d03,
     32'h000d4783,
     32'h02078863,
     32'h00000a13,
     32'h001a0a13,
     32'h014d07b3,
     32'h0007c783,
     32'hfe079ae3,
     32'h00287813,
     32'h02081a63,
     32'h001a0d93,
     32'h019a6c63,
     32'h000d8a13,
     32'h0240006f,
     32'h00000a13,
     32'hfe5ff06f,
     32'h00078d93,
     32'h02000513,
     32'hffcff0ef,
     32'h001d8793,
     32'hffbc98e3,
     32'h001c8a13,
     32'h000d0513,
     32'h869ff0ef,
     32'h001a0d13,
     32'h019a6863,
     32'h000c0a13,
     32'heb5ff06f,
     32'h00078d13,
     32'h02000513,
     32'hfccff0ef,
     32'h001d0793,
     32'hffac98e3,
     32'h000c0a13,
     32'he99ff06f,
     32'h004a0c13,
     32'h000a4503,
     32'hfb0ff0ef,
     32'h000c0a13,
     32'he85ff06f,
     32'hfa4ff0ef,
     32'he7dff06f,
     32'h00487793,
     32'h00a00693,
     32'h12079463,
     32'h00a00693,
     32'h04400793,
     32'h00f61863,
     32'h000a2703,
     32'h004a0a13,
     32'h1240006f,
     32'h000a2703,
     32'h004a0a13,
     32'h07800793,
     32'h00700893,
     32'h00f50863,
     32'h0ff8f893,
     32'h00000613,
     32'h02c0006f,
     32'h02700893,
     32'hff1ff06f,
     32'h00160c13,
     32'h018105b3,
     32'h03078793,
     32'hfef58fa3,
     32'h02d76663,
     32'h00050713,
     32'h033c0063,
     32'h000c0613,
     32'h02d777b3,
     32'h02d75533,
     32'hfcf4fce3,
     32'h00f887b3,
     32'h0ff7f793,
     32'hfcdff06f,
     32'h00f00613,
     32'h00887793,
     32'h00078c63,
     32'h01010793,
     32'h01878c33,
     32'h02d00793,
     32'hfefc0823,
     32'h00260c13,
     32'h00187793,
     32'h000b8d93,
     32'h00079463,
     32'h02000d93,
     32'h00287813,
     32'h04081463,
     32'h001c0d13,
     32'h019c6663,
     32'h01c0006f,
     32'h00078d13,
     32'h000d8513,
     32'heccff0ef,
     32'h001d0793,
     32'hffac98e3,
     32'h001c8d13,
     32'h01810c33,
     32'hfffc4503,
     32'heb4ff0ef,
     32'hfffc0c13,
     32'hff2c1ae3,
     32'h001d0c13,
     32'h019d6a63,
     32'hd7dff06f,
     32'h000c0d13,
     32'hfddff06f,
     32'h00078c13,
     32'h02000513,
     32'he8cff0ef,
     32'h001c0793,
     32'hff8c98e3,
     32'hd5dff06f,
     32'h00487793,
     32'h00098693,
     32'hee078ee3,
     32'h00098693,
     32'h004a0793,
     32'h000a2703,
     32'h04400593,
     32'h00078a13,
     32'heeb616e3,
     32'hee0754e3,
     32'h40e00733,
     32'h00886813,
     32'heddff06f,
     32'h00487793,
     32'h00200693,
     32'hea078ae3,
     32'h000a2703,
     32'h004a0a13,
     32'h00200693,
     32'hec1ff06f,
     32'h00487793,
     32'h00800693,
     32'hea0786e3,
     32'h000a2703,
     32'h004a0a13,
     32'h00800693,
     32'hea5ff06f,
     32'h04c12083,
     32'h04812403,
     32'h04412483,
     32'h04012903,
     32'h03c12983,
     32'h03812a03,
     32'h03412a83,
     32'h03012b03,
     32'h02c12b83,
     32'h02812c03,
     32'h02412c83,
     32'h02012d03,
     32'h01c12d83,
     32'h05010113,
     32'h00008067,
     32'hfc010113,
     32'h00112e23,
     32'h02b12223,
     32'h02c12423,
     32'h02d12623,
     32'h02e12823,
     32'h02f12a23,
     32'h03012c23,
     32'h03112e23,
     32'h02410593,
     32'h00b12623,
     32'hc1dff0ef,
     32'h01c12083,
     32'h04010113,
     32'h00008067,
     32'h83010113,
     32'h00112223,
     32'h00212423,
     32'h00312623,
     32'h00412823,
     32'h00512a23,
     32'h00612c23,
     32'h00712e23,
     32'h02812023,
     32'h02912223,
     32'h02a12423,
     32'h02b12623,
     32'h02c12823,
     32'h02d12a23,
     32'h02e12c23,
     32'h02f12e23,
     32'h05012023,
     32'h05112223,
     32'h05212423,
     32'h05312623,
     32'h05412823,
     32'h05512a23,
     32'h05612c23,
     32'h05712e23,
     32'h07812023,
     32'h07912223,
     32'h07a12423,
     32'h07b12623,
     32'h07c12823,
     32'h07d12a23,
     32'h07e12c23,
     32'h07f12e23,
     32'h34202573,
     32'h341025f3,
     32'h00010613,
     32'h9e1ff0ef,
     32'h00412083,
     32'h00812103,
     32'h00c12183,
     32'h01012203,
     32'h01412283,
     32'h01812303,
     32'h01c12383,
     32'h02012403,
     32'h02412483,
     32'h02812503,
     32'h02c12583,
     32'h03012603,
     32'h03412683,
     32'h03812703,
     32'h03c12783,
     32'h04012803,
     32'h04412883,
     32'h04812903,
     32'h04c12983,
     32'h05012a03,
     32'h05412a83,
     32'h05812b03,
     32'h05c12b83,
     32'h06012c03,
     32'h06412c83,
     32'h06812d03,
     32'h06c12d83,
     32'h07012e03,
     32'h07412e83,
     32'h07812f03,
     32'h07c12f83,
     32'h7d010113,
     32'h30200073,
     32'h00000093,
     32'h00008113,
     32'h00008193,
     32'h00008213,
     32'h00008293,
     32'h00008313,
     32'h00008393,
     32'h00008413,
     32'h00008493,
     32'h00008513,
     32'h00008593,
     32'h00008613,
     32'h00008693,
     32'h00008713,
     32'h00008793,
     32'h00008813,
     32'h00008893,
     32'h00008913,
     32'h00008993,
     32'h00008a13,
     32'h00008a93,
     32'h00008b13,
     32'h00008b93,
     32'h00008c13,
     32'h00008c93,
     32'h00008d13,
     32'h00008d93,
     32'h00008e13,
     32'h00008e93,
     32'h00008f13,
     32'h00008f93,
     32'h00003117,
     32'h36c10113,
     32'h00006537,
     32'h00450513,
     32'h00100593,
     32'h00b52023,
     32'h00001d17,
     32'h354d0d13,
     32'h00001d97,
     32'h364d8d93,
     32'h01bd7863,
     32'h000d2023,
     32'h004d0d13,
     32'hffbd6ce3,
     32'h00006537,
     32'h00450513,
     32'h00200593,
     32'h00b52023,
     32'h00000513,
     32'h00000593,
     32'hd3cff0ef,
     32'h0000006f,
     32'hfffff72c,
     32'hfffff78c,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7c8,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff72c,
     32'hfffff78c,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7d4,
     32'hfffff7c8,
     32'hfffffca8,
     32'hfffffb38,
     32'hfffffb54,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffcc4,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffaa8,
     32'hfffffb4c,
     32'hfffffb54,
     32'hfffffb4c,
     32'hfffffb4c,
     32'hfffffc74,
     32'h74696177,
     32'h726f6620,
     32'h726f6d20,
     32'h64252065,
     32'h63655320,
     32'h73646e6f,
     32'h000d2021,
     32'h75200a0d,
     32'h6f6e6b6e,
     32'h63206e77,
     32'h616d6d6f,
     32'h2021646e,
     32'h00000a0d,
     32'h72617453,
     32'h6f742074,
     32'h61726520,
     32'h66206573,
     32'h6873616c,
     32'h000a0d20,
     32'h72450a0d,
     32'h20657361,
     32'h706d6f43,
     32'h6574656c,
     32'h000a0d21,
     32'h3d3d0a0d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h000a0d3d,
     32'h72617473,
     32'h68742074,
     32'h70612065,
     32'h63696c70,
     32'h6f697461,
     32'h0a0d216e,
     32'h00000000,
     32'h73657250,
     32'h6e412073,
     32'h654b2079,
     32'h6f742079,
     32'h746e4920,
     32'h75727265,
     32'h42207470,
     32'h21746f6f,
     32'h00000a0d,
     32'h6d6d6f63,
     32'h20646e61,
     32'h6f727265,
     32'h0a0d2172,
     32'h00000000,
     32'h6d6d6f63,
     32'h3a646e61,
     32'h00000000,
     32'h2d2d2d2d,
     32'h2d2d2d2d,
     32'h2d2d2d2d,
     32'h6b6f6f43,
     32'h72616261,
     32'h42206172,
     32'h20746f6f,
     32'h756e654d,
     32'h2d2d2d2d,
     32'h2d2d2d2d,
     32'h2d2d2d2d,
     32'h28200a0d,
     32'h443a2944,
     32'h6c6e776f,
     32'h2064616f,
     32'h676f7250,
     32'h206d6172,
     32'h6d6f7246,
     32'h72655320,
     32'h0d6c6169,
     32'h4528200a,
     32'h72453a29,
     32'h20657361,
     32'h73616c46,
     32'h200a0d68,
     32'h3a295328,
     32'h72617453,
     32'h70412074,
     32'h000a0d70,
     32'h65637865,
     32'h6f697470,
     32'h6168206e,
     32'h656c646e,
     32'h21212172,
     32'h000a0d20,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h3d3d3d3d,
     32'h000a0d20,
     32'h544d0a0d,
     32'h3a434556,
     32'h78302020,
     32'h00000000,
     32'h454d0a0d,
     32'h203a4350,
     32'h78302020,
     32'h00000000,
     32'h434d0a0d,
     32'h45535541,
     32'h7830203a,
     32'h00000000,
     32'h544d0a0d,
     32'h3a4c4156,
     32'h78302020,
     32'h00000000,
     32'h61680a0d,
     32'h7420746c,
     32'h70206568,
     32'h65636f72,
     32'h726f7373,
     32'h00000a0d,
     32'h00000eb0,
     32'h00000ed4,
     32'h00000ee8,
     32'h00000ef4,
     32'h00000000,
     32'h00000000
    };


    // ifu read port
	always @ (*) begin
		if (rom_ce_i == `ChipDisable) begin
			rom_data_o = `ZeroWord;
		end else begin
			rom_data_o = rom_mem[rom_addr_i[`RomNumLog2+1:2]];
		end
	end

    // lsu read port
	always @ (*) begin
		if (ce_i == `ChipDisable) begin
			data_o = `ZeroWord;
	    end else if(we_i == `WriteDisable) begin
		    data_o =  rom_mem[addr_i[`RomNumLog2+1:2]];
		end else begin
			data_o = `ZeroWord;
		end
	end

/*
    // Task for loading 'rom_mem' with SystemVerilog system task $readmemh()
    export "DPI-C" task simutil_romload;

    task simutil_romload;
        input string file;
        $readmemh(file, rom_mem);
    endtask

    // Function for setting a specific element in |rom_mem|
    // Returns 1 (true) for success, 0 (false) for errors.
    export "DPI-C" function simutil_set_rom;

    function int simutil_set_rom(input int index, input bit [`InstBus] val);
        if (index >= `RomNum) begin
            return 0;
        end
        rom_mem[index] = val;
        return 1;
    endfunction

    // Function for getting a specific element in |rom_mem|
    export "DPI-C" function simutil_get_rom;

    function int simutil_get_rom(input int index, output bit [31:0] val);
        if (index >= `RomNum) begin
          return 0;
        end

        val = 0;
        val = rom_mem[index];
        return 1;
    endfunction
*/

endmodule
